-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Oct 20 17:35:34 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Motor_c_ADCs IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Der_Cerca : IN STD_LOGIC := '0';
        Izq_Cerca : IN STD_LOGIC := '0';
        MD : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        MI : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END Motor_c_ADCs;

ARCHITECTURE BEHAVIOR OF Motor_c_ADCs IS
    TYPE type_fstate IS (Avanza,Izquierda_cerca,Derecha_cerca);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Der_Cerca,Izq_Cerca)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Avanza;
            MD <= "00";
            MI <= "00";
        ELSE
            MD <= "00";
            MI <= "00";
            CASE fstate IS
                WHEN Avanza =>
                    IF (((Der_Cerca = '0') AND (Izq_Cerca = '0'))) THEN
                        reg_fstate <= Avanza;
                    ELSIF (((Der_Cerca = '1') AND (Izq_Cerca = '0'))) THEN
                        reg_fstate <= Derecha_cerca;
                    ELSIF ((Izq_Cerca = '1')) THEN
                        reg_fstate <= Izquierda_cerca;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Avanza;
                    END IF;

                    MD <= "01";

                    MI <= "01";
                WHEN Izquierda_cerca =>
                    IF (((Izq_Cerca = '0') AND (Der_Cerca = '1'))) THEN
                        reg_fstate <= Derecha_cerca;
                    ELSIF (((Izq_Cerca = '0') AND (Der_Cerca = '0'))) THEN
                        reg_fstate <= Avanza;
                    ELSIF ((Izq_Cerca = '1')) THEN
                        reg_fstate <= Izquierda_cerca;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Izquierda_cerca;
                    END IF;

                    MD <= "10";

                    MI <= "01";
                WHEN Derecha_cerca =>
                    IF (((Izq_Cerca = '1') AND (Der_Cerca = '0'))) THEN
                        reg_fstate <= Izquierda_cerca;
                    ELSIF (((Der_Cerca = '0') AND (Izq_Cerca = '0'))) THEN
                        reg_fstate <= Avanza;
                    ELSIF ((Der_Cerca = '1')) THEN
                        reg_fstate <= Derecha_cerca;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Derecha_cerca;
                    END IF;

                    MD <= "01";

                    MI <= "10";
                WHEN OTHERS => 
                    MD <= "XX";
                    MI <= "XX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
